module json

pub fn decode(typ voidptr, s string) ?voidptr {
	// compiler implementation
	return 0
}

pub fn encode(x voidptr) string {
	// compiler implementation
	return ''
}
