module builtin

pub struct array {
pub:
	len int
}
