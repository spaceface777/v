// Copyright (c) 2019-2020 Alexander Medvednikov. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module pref

pub enum OS {
	_auto // Reserved so .mac cannot be misunderstood as auto
	ios
	mac
	linux
	windows
	freebsd
	openbsd
	netbsd
	dragonfly
	js // TODO
	android
	solaris
	haiku
}

// Helper function to convert string names to OS enum
pub fn os_from_string(os_str string) ?OS {
	match os_str {
		'linux' {
			return .linux
		}
		'windows' {
			return .windows
		}
		'ios' {
			return .ios
		}
		'mac' {
			return .mac
		}
		'macos' {
			return .mac
		}
		'freebsd' {
			return .freebsd
		}
		'openbsd' {
			return .openbsd
		}
		'netbsd' {
			return .netbsd
		}
		'dragonfly' {
			return .dragonfly
		}
		'js' {
			return .js
		}
		'solaris' {
			return .solaris
		}
		'android' {
			return .android
		}
		'haiku' {
			return .haiku
		}
		'linux_or_macos' {
			return .linux
		}
		'' {
			return ._auto
		}
		else {
			return error('bad OS $os_str')
		}
	}
}

pub fn (o OS) str() string {
	match o {
		._auto {
			return 'RESERVED: AUTO'
		}
		.ios {
			return 'iOS'
		}
		.mac {
			return 'MacOS'
		}
		.linux {
			return 'Linux'
		}
		.windows {
			return 'Windows'
		}
		.freebsd {
			return 'FreeBSD'
		}
		.openbsd {
			return 'OpenBSD'
		}
		.netbsd {
			return 'NetBSD'
		}
		.dragonfly {
			return 'Dragonfly'
		}
		.js {
			return 'JavaScript'
		}
		.android {
			return 'Android'
		}
		.solaris {
			return 'Solaris'
		}
		.haiku {
			return 'Haiku'
		}
	}
}

pub fn get_host_os() OS {
	$if linux           { return linux }
	$else $if ios       { return ios }
	$else $if macos     { return mac }
	$else $if windows   { return windows }
	$else $if freebsd   { return freebsd }
	$else $if openbsd   { return openbsd }
	$else $if netbsd    { return netbsd }
	$else $if dragonfly { return dragonfly }
	$else $if solaris   { return solaris }
	$else $if haiku     { return .haiku }
	panic('unknown host OS')
}
